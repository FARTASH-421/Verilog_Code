// module LeftControl (
//     input rest, clk,
//     input [3:0] F
//     input [3:0] Up, Down, 
//     input [3:0] S,

//     output [2:0] AC,
//     output [4:0] DISP,
//     output open
// );



// always@(posedge clk or posedge rst )
// begin
// 	if (rst)begin
//         AC = 0;
//         DISP = 0;
//         open = 0;
// 	end
// 	else begin
//     if()

//     end
// end
    
// endmodule